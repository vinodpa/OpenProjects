

module tb_avalon ();

endmodule